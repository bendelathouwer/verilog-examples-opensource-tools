`timescale 1ns/1ps
module clockdevider_tb(output wire o_led);



endmodule