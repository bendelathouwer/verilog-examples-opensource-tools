`timescale 1ns/100ps
module buttoncounter_TB;
reg button;
reg clk
wire [6:0] display;
buttoncounter u1 
(
        
)
endmodule